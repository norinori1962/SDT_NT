************************************************
* Export Spice: 
* Library Name: sim_tsuda
* Top Cell Name: git_test
* Netlisted on: Fri Jun 24 16:43:24 2016
*				 JEDAT Inc.
************************************************

************************************************
* DUT: sim_tsuda/git_test/schematic
************************************************


************************************************
*sim_tsuda/git_test
************************************************

*.SUBCKT git_test IN OUT 
r000 IN OUT 2K

*----------------------------------------------*
*      Cross Reference List for node No.       *
*----------------------------------------------*
*          name                    No.


*.ENDS git_test


************************************************
* .PARAM
************************************************
.END
